*
**********************************************************
*
* PSSI2021SAY
*
* NXP Semiconductors
*
* Constant current source
* output current = max 50mA
* supply voltage = max 75V 
*
*
*
*
*
* Package pinning does not match Spice model pinning.
* Package: SOT 353
*  
* Package Pin 1: not connected   4: external resistor
* Package Pin 2: output current  5: supply voltage
* Package Pin 3: GND
*
* 
*
* Simulator: Spice 2
*
**********************************************************
*#
.SUBCKT PSSI2021SAY 1 2 3 4
*
Q1 1 22 3 MAIN
D1 4 44 DIODE1
D2 44 22 DIODE2
RD2 44 22 5E+09
Rbase 2 22 3.35E+04
Rint 3 4 5.28E+04
*
.MODEL MAIN PNP
+ IS = 4.512E-14
+ NF = 1.004
+ ISE = 1E-25
+ NE = 0.9237
+ BF = 120
+ IKF = 1.1
+ VAF = 104
+ NR = 1.002
+ ISC = 1.465E-11
+ NC = 1.599
+ BR = 16.5
+ IKR = 5E+04
+ VAR = 12.7
+ RB = 27
+ IRB = 0.00074
+ RBM = 1.595
+ RE = 0.1
+ RC = 0.23
+ XTB = 0
+ EG = 1.11
+ XTI = 3
+ CJE = 0
+ VJE = 0.75
+ MJE = 0.333
+ TF = 2E-30
+ XTF = 0
+ VTF = 1000
+ ITF = 0
+ PTF = 0
+ CJC = 0
+ VJC = 0.75
+ MJC = 0.333
+ XCJC = 1
+ TR = 1E-32
+ CJS = 0
+ VJS = 0.75
+ MJS = 0.333
+ FC = 0.78
.MODEL DIODE1 D
+ IS = 1.673E-14
+ N = 1.089
+ BV = 1000
+ IBV = 0.001
+ RS = 0.7739
+ CJO = 0
+ VJ = 1
+ M = 0.5
+ FC = 0
+ TT = 0
+ EG = 1.11
+ XTI = 3
.MODEL DIODE2 D
+ IS = 1.12E-14
+ N = 1.076
+ BV = 1000
+ IBV = 0.001
+ RS = 0.8848
+ CJO = 0
+ VJ 1
+ M = 0.5
+ FC = 0
+ TT = 0
+ EG = 1.11
+ XTI = 3
.ENDS