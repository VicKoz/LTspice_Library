* ADA4850 SPICE Macro-model        
* Description: Amplifier
* Generic Desc: LC Voltage Feedback RR Dual w/Disable
* Developed by:
* Revision History: 08/10/2012 - Updated to new header style
*
* Copyright 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model 
* indicates your acceptance of the terms and provisions in the License Statement.
* 
* BEGIN Notes:
*
* Not Modeled:
*    
* Parameters modeled include: 
* END Notes
*
* Node assignments

.SUBCKT ADA4850 NINV INV VCC VEE OUT  
***************************************
* Analog Devices ADA4850
* 2005.05.25 v1.1
****************************************
*  Features included in model
* 1. Open loop gain and phase
* 2. Output voltage and current
* 3. Input Common mode range
* 4. Input Bias current
* 5. Input voltage and current noise
* 6. Slew rate
* 7. Output current reflected in Vs supplies
* 8. Transient Response
* 9. Frequency Response
***************************************
Q_Q1         V5 92 7 NPN 
Q_Q2         V6 INV 8 NPN 
R_RC1         VCC_INT V5 RCOLD 101.034
R_RC2         VCC_INT V6 RCOLD 101.034
R_RE1         7 4 RCOLD 100
R_RE2         8 4 RCOLD 100
I_I1         4 VEE_INT DC .05  
E_EOS         NINV 9 POLY(1) CMRR_V 100 0.0 1
E_ENIN         92 9 36 0 2.5e-7
G_G8         100 CMRR_V CMRRP2 100 .01
G_G7         100 CMRRP2 CMRRP1 100 .01
G_G6         100 CMRRP1 30 100 .01
R_RCM         31 100 RCOLD 1E2
R_RCM1         NINV VINMID RCOLD 1000MEG
R_RCM2         VINMID INV RCOLD 1000MEG
R_RCM2a         CMRRP1 100 RCOLD 100
C_CCM2a         100 CMRRP1  2.6526e-11  
R_RCM3         CMRRP2 100 RCOLD 100
C_CCM3         100 CMRRP2  1.9894e-11  
R_RCM4         CMRR_V 100 RCOLD 100
C_CCM4         100 CMRR_V  1.9894e-12  
L_LCM         31 30  2.274e-3  
R_RP1         10 100 RCOLD 100
C_CP1         100 10  8.07e-6  
R_RP2         N10305 100 RCOLD 100
C_CP2         100 N10305  1.326e-11  
R_RP3         MAINP2 100 RCOLD 100
C_CP3         100 100  1.0610e-12  
V_VN         VEEVNBAT VEE_INT .505
V_VN1         0 35 2Vdc
D_DN5         96 97 DIN 
V_V1         VCC_INT N129837 2.7
D_DN1         35 36 DEN 
D_DN3         93 94 DIN 
V_VN2         37 0 2Vdc
D_DN2         36 37 DEN
V_VN3         0 93 2
D_DN4         94 95 DIN 
V_VN4         95 0 2
G_GN1         0 NINV 94 0 2.15e-9
V_VN5         0 96 2
D_DN6         97 98 DIN 
V_VN6         98 0 2
R_R3         ISUPP1 0 RCOLD 10meg
D_D_VEEclamp         VEEVNBAT 10 DN 
D_D_VCCclamp         10 VCCVPBAT DP 
D_D7         ISUPP2 0 DZ 
C_C1         100 81  4p  
E_E5         VEE_INT 0 VEE 0 1
G_G2         100 N10305 10 100 1e-2
G_G1         100 10 N06761 100 7.1
D_D8         VCC ISUPP1 DNOM 
G_GV         100 N06761 V6 V5 .001
E_E6         103 VEE_INT VALUE { (V(VCC_INT)-V(VEE_INT))/2 }
V_VP         VCC_INT VCCVPBAT .499
G_G3a         100 MAINP2 N10305 100 1e-2
D_D9         ISUPP2 VEE DNOM 
E_E4         VCC_INT 0 VCC 0 1
R_R4         0 ISUPP2 RCOLD 10meg
D_D5         INV N129837 DP 
G_G5         100 30 VINMID 100 3.162e-8
D_DZ2         100 16 DLIM 
D_DZ1         N06761 16 DLIM 
G_G10         0 INV 97 0 2.15e-9
G_G3         ISUPP1 0 80 81 .02
G_G4         0 ISUPP2 80 81 -.02
I_IQP         ISUPP1 0 DC 2.5m  
I_IQM         0 ISUPP2 DC 2.5m  
D_D6         0 ISUPP1 DZ 
E_E1         100 0 103 0 1
E_EBUF         80 100 MAINP2 100 1
L_Lout         OUT 81  60n  
R_Rout         80 81 RCOLD 50
R_RV         N06761 100 RCOLD 500k
.MODEL DLIM D(IS=1E-15 BV=1010)
.MODEL DEN  D(IS=1E-8 RS=1 KF=1E-15 AF=1)
.MODEL DIN  D(IS=.75E-12 RS=100 KF=3e-15 AF=1)
.MODEL	DNOM	D(IS=1E-15 T_ABS=-100)
.MODEL	DZ	D(IS=1E-15 BV=50 T_ABS=-100)
.MODEL  RCOLD	RES T_ABS=-273
.MODEL 	DILIM	D(IS=1E-15)
.MODEL NPN  NPN(BF=1.47e4)
.MODEL	DP	D(IS=5E-10 BV=700 )
.MODEL	DN	D(IS=5E-10 BV=700 )
.ENDS




