* AD8638 SPICE Macro-model Typical Values
* Description: Amplifier
* Generic Desc: 5/16V, CMOS, OP, Zero Drift, S SPLY, 1X
* Developed by: HH/ADISJ
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (11/2007)
* Copyright 2007, 2012 by Analog Devices
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement.  Use of this model
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*    
* Parameters modeled include: 
*
* END Notes
*
* Node Assignments
*                       noninverting input
*                       |   inverting input
*                       |   |    positive supply
*                       |   |    |   negative supply
*                       |   |    |   |   output
*                       |   |    |   |   |
*                       |   |    |   |   |
.SUBCKT AD8638          1   2   99  50  45
*
* INPUT STAGE
*
M1  14  7  8  8 PIX L=1E-6 W=2.092E-05
M2  16  2  8  8 PIX L=1E-6 W=2.092E-05
RC5 14 50 1.200E+04
RC6 16 50 1.200E+04
C1  141 16 1.300E-12
RC56 14 141 2.0E-04
I1  99  8 5.000E-05
V1  99  9 2.001E+00
D1   8  9 DX
EOS  7  1 POLY(4) (22,98) (73,98) (83,98) (70,98) 3.00E-06 1 1 1.275 1
IOS  1  2 5.00E-12
*
* CMRR=140dB, POLE AT 12.5 Hz
*
E1  21 98 POLY(2) (1,98) (2,98) 0 2.066E-02 2.066E-02
R10 21 22 1.315E+04
R20 22 98 3.183E-02
C10 21 22 1.000E-06
*
* PSRR=143dB, POLE AT 0.1 Hz
*
EPSY 72 98 POLY(1) (99,50) -26.1395E+00 1.67337E+00
RPS3 72 73 1.224E+06
RPS4 73 98 5.305E-02
CPS3 72 73 1.00E-06
*
* VOLTAGE NOISE REFERENCE OF 60nV/rt(Hz)
*
VN1 80 98 0
RN1 80 98  80.0E-06
*
HN  81 98 VN1 220E+00
RNHH1 81 183 5.3
CHH1 183 98 1uF
*
CHH2 183 184 2.7E-07
RNHH2 184 98 10
*
RNHH3 184 83 129k
CHH3 83 98 2.41E-10
*
* FLICKER NOISE CORNER = 0.0001 Hz
*
D5  69 98 DNOISE
VSN 69 98 DC 0.6551
H1  70 98 POLY(1) VSN 1.00E-03 1.00E+00
RN  70 98 1
*
* INTERNAL VOLTAGE REFERENCE
*
EREF 98  0 POLY(2) (99,0) (50,0) 0 0.5 0.5
GSY  99 50 POLY(1) (99,50) 0.7151E-03 8.763E-06
EVP  97 98 POLY(1) (99,50) 0 0.5E-09
EVN  51 98 POLY(1) (50,99) 0 0.5E-09
*
* GAIN STAGE
*
G1 98 130 POLY(1) (14,16)  0 2.054E-01
RG1 130 30 1
R1 30 98 1.00E+06
CR1 30 98 1.00E-15
V3 32 30 -0.429E+00
V4 30 33 -1.560E+00
*
EZ (145 0) POLY(1) (45 0) 0 1
REZ 145 0 10Meg
*
CF 145 31 5.950E-08
RZ 30 31 1.00E-01
D3 32 97 DX
D4 51 33 DX
*
* OUTPUT STAGE
*
M5  45 46 99 99 POX L=1E-6 W=1.455E-04
M6  45 47 50 50 NOX L=1E-6 W=1.875E-04
EG1 99 46 POLY(1) (98,30) 5.626E-01 1
EG2 47 50 POLY(1) (30,98) 4.966E-01 1
*
* MODELS
*
.MODEL POX PMOS (LEVEL=2,KP=5.00E-05,VTO=-0.4,LAMBDA=0.05,RD=0.5)
.MODEL NOX NMOS (LEVEL=2,KP=11.00E-05,VTO=+0.4,LAMBDA=0.04,RD=0.7)
.MODEL PIX PMOS (LEVEL=2,KP=5.00E-05,VTO=-6.00E-01,LAMBDA=0.02)
.MODEL DX D(IS=1E-14,RS=5)
.MODEL DNOISE D(IS=1E-14,RS=0,KF=2.50E-20)
*
*
.ENDS AD8638
*
*$




