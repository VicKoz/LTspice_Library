* ADA4930 SPICE Macro-model
* Description: Amplifier
* Generic Desc: UltraLow Dist Low Vltg ADC Driver
* Developed by: CK
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (07/2011)
* Copyright 2006, 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*     distortion is not characterized
*     cmrr is not characterized in this version.
*
* Parameters modeled include:
*     closed loop gain and phase vs bandwidth
*     output current and voltage limiting
*     offset voltage (is  non-static, will  vary with gain)
*     ibias (again, is static, will not vary with vcm)
*     slew rate and step response performance
*     (slew rate is based on 10-90% of step response)
*     current on output will be reflected to the supplies 
*     Vocm is varable and include input typical offset
*     Voltage Noise in also included.
*
* END Notes:
*
* Node assignments
*               FD output negative
*                | FD output positive
* 		 | |  non-inverting input
*		 | |  | inverting input
*		 | |  |  |  positive supply
*		 | |  |  |  |  negative supply
*		 | |  |  |  |  |  output positive
*		 | |  |  |  |  |  |   output negative
*		 | |  |  |  |  |  |   |   vocm input
*		 | |  |  |  |  |  |   |   |
.SUBCKT ADA4930 9b 3b 3a 9 99 50 71b 71  110

*** positive input left side ***

I 99 5 8E-4
Q1 50 2 5 QX
vos 3a 2 -1.95E-3

*** RAIL CLIPING ***

Dlim+ 75a 14b Dx
Vlim+ 99 14b 2.28
Dlim 14c 75a Dx
Vlim 14c  50 1.08
Dlim- 13b 76a DX
Vlim- 13b 50 1.08
Dlim-B 76a 13C Dx
Vlim-B 99 13C 2.28

*** VOCM INPUT RAIL CLIPING ***

DOCMa 100 100a dx
VOCMa 99 100a 2.81
DOCMb 100b 100 DX
VOCMb 100b 50 1.35

*** negative input right side ***

I1 99 6 8E-4
Q2 50 9 6 QX

*** Input capacitance/impedance ***

Cin 3a 9 0.6p

*** pole, zero pole stage ***

G1 13 14 5 6 5E-3
c1 14 13 80f
c2 98 13 700f
c3 98 14 700f
r11 98 13 RX1 250K 
r12 98 14 RX1 250K 

*** pole zero stage( POSITIVE SIDE) ***

gp1 0 75 14 98 1
RP1 75 0 RX2 1
CP1 0 75 0.1p

*** pole zero stage( NEGATIVE SIDE) ***

gp2 0 76 13 98 1
RP2 76 0 RX2 1
CP2 0 76 0.1pf

*** output stage Negative side ***

D17 76 84 DX
VO1  84 70 .177V
VO2  70 85 .177V
D16 85 76  DX
G30 70 99c 99 76  91E-3
G31 98c 70 76 50  91E-3
RO30 70 99c RX2 11
RO31 98c 70 RX2 11 
VIOUT1 99 99c 0
VIOUT2 98c 50 0
VIOUT3 70 71 0

*** Output Stage Positive side ***

D17b 75 84b DX
VO1b  84b 70b .177V
VO2b  70b 85b .177V
D16b 85b 75  DX
G30b 70b 99d 99 75  91E-3
G31b 98d 70b 75 50  91E-3
RO30b 70b 99d RX2 11
RO31b 98d 70b RX2 11 
VIOUTB1 99 99d 0
VIOUTB2 98d 50 0
VIOUTB3 70b 71b 0

*** VOCM STAGE ***

Gocm_a 0 75 100 0 1
Gocm_b 0 76 100 0 1
Rocm1 110 99 20K 
Rocm2 50 110 20K 

Voffset 100 110 -10E-3

*** CURRENT MIRROR TO SUPPLIES POSITVIE SIDE ***

FO1 0 99 poly(2) VIOUT1 VI1 -17.503E-3 1 -1
FO2 0 50 poly(2) VIOUT2 VI2 -17.503E-3 1 -1
FO3 0 400 VIOUT1 1
VI1 401 0 0
VI2 0 402 0
DM1 400 401 DX
DM2 402 400 DX 

*** CURRENT MIRROR TO SUPPLIES NEGATIVE SIDE ***

FO1B 0 99 poly(2) VIOUTB1 VIB1 -16E-3 1 -1
FO2B 0 50 poly(2) VIOUTB2 VIB2 -16E-3 1 -1
FO3B 0 400B VIOUTB1 1
VIB1 401B 0 0
VIB2 0 402B 0
DMB1 400B 401B DX
DMB2 402B 400B DX

*** Reference Stage ***

Eref 98 0 poly(2) 99 0 50 0 0 0.5 0.5

*** Feadback output ***

Vfd+ 3b 71b 0
Vfd- 9b 71  0

*** Buffer Stage ***

Vbf1 76 76a 0
Vbf2 75 75a 0

*** Models ***

.MODEL QX PNP (BF=228 Is=1E-15 KF=1E-12 AF=1.0)
.MODEL RX1 Res(T_abs=-0)
.MODEL RX2 Res(T_abs=-0)
*.MODEL RX3 Res(T_abs=-0)
.MODEL DX D(IS=1E-14)
*.MODEL DEN D(IS=1E-9 RS=0.004 KF=7E-10 AF=1)
.ENDS
;$SpiceType=AMBIGUOUS
*$




