* OPA191 Spice simulation model
*
* Copyright 2015 by Texas Instruments Corporation
*
* OPA191 Rev A, by Tim Green; December 10, 2015
*
* This macromodel has been optimized to model the AC, DC, noise,
* and transient response performance within the device data sheet
* specified limits. Correct operation of this macromodel has been
* verified on DesignSoft TINA Version 7.0.80.224 SF and Penzar 
* TopSPICE 8, version 8.39. For help with other analog simulation
* software, please consult the software supplier.
*
* BEGIN MODEL OPA191
*
* GREEN-LIS MACRO-MODEL SIMULATED FEATURES:
*
* OPEN LOOP GAIN AND PHASE VS FREQUENCY WITH RL AND CL EFFECTS
* INPUT COMMON MODE REJECTION WITH FREQUENCY
* POWER SUPPLY REJECTION WITH FREQUENCY
* INPUT IMPEDANCE VS FREQUENCY 
* OUTPUT IMPEDANCE VS FREQUENCY 
* INPUT VOLTAGE NOISE VS FREQUENCY
* INPUT CURRENT NOISE VS FREQUENCY 
* OUTPUT VOLTAGE SWING VS OUTPUT CURRENT
* SHORT-CIRCUIT OUTPUT CURRENT
* QUIESCENT CURRENT VS SUPPLY VOLTAGE
* SETTLING TIME VS CAPACITIVE LOAD
* SLEW RATE
* SMALL SIGNAL OVERSHOOT VS CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME
* INPUT BIAS CURRENT
* INPUT VOLTAGE OFFSET
* INPUT COMMON MODE RANGE
* OUTPUT CURRENT COMING THROUGH THE SUPPLY RAILS
*
.SUBCKT OPA191 +IN -IN V+ V- Vout
V6          V- 38 -200M
V5          37 V+ -200M
V1          71 Vee_B -100M
VscNeg      MID 73 1
V3          MID 76 300
V2          77 MID 300
V12         MID 83 64.2
V8          84 MID 64.2
V7          85 Vcc_B 100M
IS2         +PSR V- 5P
Vos         -CMR 36 -30.9656U
VscPos      75 MID 1
VoldPos     74 MID 7.6
VoldNeg     MID 72 2.8
Iq          V+ V- 140U
IS3         80 V- 3P
XU17        33 MID 34 MID VCVS_LIMIT_0
XVn11       35 36 VNSE_0
XIn11       36 -IN_F FEMT_0
R8          +CMR -PSR 1M 
XD1         Vout V+ D_D_0
XD2         V- Vout D_D_0
R30         +CMR -CMR 1G 
R1          +PSR -PSR 1G 
XT1         37 -CMR 37 JFET_TG_0
XT2         -CMR 38 -CMR JFET_TG_0
XT3         37 -IN_F 37 JFET_TG_0
XT4         -IN_F 38 -IN_F JFET_TG_0
GVCCS22     39 40 39 40  1.01U
GVCCS21     41 42 41 42  1.01U
GVCCS20     43 44 43 44  1.01U
GVCCS19     MID 45 MID 45  180.65U
GVCCS18     MID 46 MID 46  22.08
GVCCS17     47 40 47 40  100U
GVCCS16     48 45 48 45  100U
GVCCS14     49 46 49 46  100U
EVCVS12     39 MID 45 MID  2.806452
C19         48 45 25.67015P 
EVCVS11     48 MID 46 MID  220.8122K
R15         MID 40 1G 
C18         MID 47 32.54702F 
C14         49 46 2.019733U 
EVCVS9      49 MID Vee_B MID  1U
GVCCS13     MID 50 MID 50  180.65U
GVCCS12     MID 51 MID 51  22.08
GVCCS11     52 42 52 42  100U
GVCCS10     53 50 53 50  100U
GVCCS9      54 51 54 51  100U
EVCVS10     41 MID 50 MID  2.806452
C17         53 50 25.67015P 
EVCVS8      53 MID 51 MID  220.8122K
R12         MID 42 1G 
C16         MID 52 32.54702F 
C15         54 51 2.019733U 
EVCVS6      54 MID Vcc_B MID  1U
GVCCS8      44 55 44 55  100U
GVCCS4      56 MID 56 MID  4.1694
GVCCS3      57 56 57 56  100U
EVCVS5      +CMR -CMR 44 MID  1
EVCVS4      43 MID 56 MID  131.7552M
R29         MID 44 1G 
C8          MID 55 44.70644F 
C3          57 56 1.070309U 
EVCVS2      57 MID -CMR MID  1
SW1         58 59 OLD_SW MID  S_VSWITCH_1
C13         Zo_out MID  3.70000000000000E-0016 
R26         MID 60 1G 
R25         61 60 20.71429K 
C11         MID 62 740.2555F 
R24         62 60 10K 
EVCVS1      61 MID 63 MID  1
C9          64 65 36.25397P 
R23         MID 65 3.348589K 
R22         64 65 10K 
EStage_1    64 MID 58 MID  2.4
RC2         MID 63 1G 
C4          66 33 636.6198F 
R11         MID 33 114.9425 
R10         66 33 10K 
R9          67 63 20.71429K 
C2          MID 68 740.2555F 
R7          68 63 10K 
EStage_3    66 MID 60 MID  1
C1          59 58 53.05165U 
R6          MID 58 7.142857K 
R5          59 58 10K 
EStage_2    67 MID 65 MID  3.986333
EDC         59 MID Zo_in Zo_out  90
Rdummy      MID Zo_out 33K 
Rx          34 Zo_out 333K 
XR109       Vsense MID RNOISE_FREE_0
XR109_2     Jaol MID RNOISE_FREE_0
C5          MID 69 4P IC=0 
R2          Vimon 69 100 
C10         MID 70 4P 
R21         Vimon 70 100 
XU7         MID OVLD- 72 Vclp 73 SC- OVLD_THRES_0
XU2         MID OVLD+ 74 Vclp 75 SC+ OVLD_THRES_0
XU16        MID OLD_SW OL+ OL- OL_CNTL_0
XU15        70 MID V- MID VCCS_LIMIT_0
XU14        70 MID V+ MID VCCS_LIMIT_1
XU3         OVLD+ OVLD- Vsense MID OL+ OL- CLMP_AMP_0
XU1         OL+ OL- Over_clamp MID VCCS_LIMIT_2
XU13        77 76 Over_clamp MID 78 79 CLMP_AMP_0
XU12        78 79 Over_clamp MID VCCS_LIMIT_2
R4          -IN_F 80 1M 
XU11        VCC_CLP VEE_CLP Vout MID 81 82 CLMP_AMP_0
XU10        81 82 CLAW_clamp MID VCCS_LIMIT_3
XU9         84 83 69 MID SC+ SC- CLMP_AMP_0
XU8         SC+ SC- CL_clamp MID VCCS_LIMIT_3
XVcm        +PSR 86 85 71 VCVS_EXT_LIMIT_0
EVCVS7      +PSR -PSR 42 40  1
R3          0 87 1G 
GVCCS7      87 Vee_B 87 Vee_B  1U
GVCCS2      87 Vcc_B 87 Vcc_B  1U
VCCVS1_in   Zo_out Vout
HCCVS1      Vimon MID VCCVS1_in   1K
C7          -IN_F 35 1.6P IC=-504.1045803864U 
Ccmp        35 MID 6.4P IC=1.000702095 
Ccmm        MID -IN_F 6.4P IC=-1.0001979904 
XR109_3     CLAW_clamp MID RNOISE_FREE_0
XU5         Vimon MID V+ VCC_CLP VCVS_LIMIT_1
XU6         MID Vimon VEE_CLP V- VCVS_LIMIT_2
C23         MID Vclp 4P IC=0 
R13         Zo_in Vclp 100 
GVCCS1      MID CLAW_clamp Jaol MID  1M
XU26        86 80 MID 88 VCCS_LIMIT_4
XU4         88 MID 0 Over_clamp VCCS_LIMIT_5
XR109_4     CL_clamp MID RNOISE_FREE_0
GVCCS15     MID CL_clamp CLAW_clamp MID  1M
R20         +IN 35 10M 
R18         -IN -IN_F 10M 
GVCCS6      MID Jaol Vsense MID  1M
C6          87 0 1 IC=0 
XR104       Over_clamp 0 RNOISE_FREE_1
XR103       MID 88 RNOISE_FREE_1
EVCVS34     MID 0 87 0  1
EVCVS29     Vcc_B 0 V+ 0  1
EVCVS28     Vee_B 0 V- 0  1
GVCCS5      MID Vsense Over_clamp MID  1M
Ccc         Over_clamp 0 784.5N IC=1.0032648632 
EVCVS3      Zo_in MID CL_clamp MID  1
.MODEL S_VSWITCH_1 VSWITCH (RON=100U ROFF=1T VON=900M VOFF=100M)
.ENDS


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_0  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 88
.PARAM VPOS = 21.8K
.PARAM VNEG = -21.8K
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VNEG,VPOS)}
.ENDS VCVS_LIMIT_0 


* BEGIN PROG NSE NANO VOLT/RT-HZ
.SUBCKT VNSE_0  1 2
* BEGIN SETUP OF NOISE GEN - NANOVOLT/RT-HZ
* INPUT THREE VARIABLES
* SET UP VNSE 1/F
* NV/RHZ AT 1/F FREQ
.PARAM NLF=48
* FREQ FOR 1/F VAL
.PARAM FLW=100
* SET UP VNSE FB
* NV/RHZ FLATBAND
.PARAM NVR=19
* END USER INPUT
* START CALC VALS
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
* END CALC VALS
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS
* END PROG NSE NANOV/RT-HZ


* BEGIN PROG NSE FEMTO AMP/RT-HZ 
.SUBCKT FEMT_0  1 2
* BEGIN SETUP OF NOISE GEN - FEMPTOAMPS/RT-HZ
* INPUT THREE VARIABLES
* SET UP INSE 1/F
* FA/RHZ AT 1/F FREQ
.PARAM NLFF=1.5
* FREQ FOR 1/F VAL
.PARAM FLWF=1E-3
* SET UP INSE FB
* FA/RHZ FLATBAND
.PARAM NVRF=1.5
* END USER INPUT
* START CALC VALS
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
* END CALC VALS
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS
* END PROG NSE FEMTO AMP/RT-HZ


.LIB "C:\Program Files (x86)\Tina Industrial 9.3\SPICELIB\ICDEVS.LIB"
*
* CONNECTIONS:   A
*                |    C
*                |    |
.SUBCKT D_D_0       1    2
D1 1 2  DCO
.MODEL DCO D RS=20 CJO=0.1E-12 TT=1E-8
.ENDS D_D_0 


*JFET FOR CLAMP DIODES IN GREEN-LIS OP AMP MACRO-MODEL
.SUBCKT JFET_TG_0  D G S
JIDEAL D G S NJFET
.MODEL NJFET NJF RD=10 RS=10 IS=1E-18
.ENDS JFET_TG_0 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_0  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E3
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_0 


* OVERLOAD THRESHOLD CONTROL FOR GL MACRO MODEL
.SUBCKT OVLD_THRES_0  1   2    3    4    5  6 
*PINS             COM OVLD VOLD VCLP VSC SC
ESW 2 1 VALUE = {IF( (V(6,1)>100M),(V(4,1)+V(5,1)), (V(4,1)+V(3,1)) )}
.ENDS OVLD_THRES_0 


* CLAMP AMP FOR CONTROL OF EXTERNAL VCCS
.SUBCKT OL_CNTL_0  1   2  3    4 
*PINS          COM SW OLD+ OLD-
ESW 2 1 VALUE = {IF((V(3,1)>10U | V(4,1)>10U),1,0)}
.ENDS OL_CNTL_0 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_0  VC+ VC- IOUT+ IOUT-
*              
.PARAM GAIN = 1M
*.PARAM IPOS = 50M
*.PARAM INEG = 0
G1 IOUT+ IOUT- VALUE={IF( (V(VC+,VC-)>=0),0,GAIN*V(VC+,VC-) )}
*G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
*ESW 2 1 VALUE = {IF( (V(6,1)>100M),(V(4,1)+V(5,1)), (V(4,1)+V(3,1)) )}
.ENDS VCCS_LIMIT_0 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_1  VC+ VC- IOUT+ IOUT-
*              
.PARAM GAIN = 1M
*.PARAM IPOS = 50M
*.PARAM INEG = 0
G1 IOUT+ IOUT- VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
*G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
*ESW 2 1 VALUE = {IF( (V(6,1)>100M),(V(4,1)+V(5,1)), (V(4,1)+V(3,1)) )}
.ENDS VCCS_LIMIT_1 


* CLAMP AMP FOR CONTROL OF EXTERNAL VCCS
.SUBCKT CLMP_AMP_0  VC+ VC- VIN COM VO+ VO-
*  TERMINALS     CLAMP V+  CLAMP V-  VIN  VOUT+  VOUT-
.PARAM G=100
EVO+ VO+ COM VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
EVO- VO- COM VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS CLMP_AMP_0 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_2  VC+ VC- IOUT+ IOUT-
*              
.PARAM GAIN = 1
.PARAM IPOS = 100
.PARAM INEG = -100
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS VCCS_LIMIT_2 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_3  VC+ VC- IOUT+ IOUT-
*              
.PARAM GAIN = 1M
.PARAM IPOS = 400M
.PARAM INEG = -400M
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS VCCS_LIMIT_3 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_EXT_LIMIT_0  VIN VOUT VP+ VP-
*              
.PARAM GAIN = 1
E1 VOUT 0 VALUE={LIMIT(GAIN*V(VIN,0),V(VP+,0),V(VP-,0))}
.ENDS VCVS_EXT_LIMIT_0 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_1  VC+ VC- VOUT+ VOUT-
*              
E1 VOUT+ VOUT- TABLE {ABS(V(VC+,VC-))} = 
+(0, 5E-3)
+(40, 1.8)
+(62, 3.37)
+(80, 6.42)
.ENDS VCVS_LIMIT_1 



*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_2  VC+ VC- VOUT+ VOUT-
*              
E1 VOUT+ VOUT- TABLE {ABS(V(VC+,VC-))} = 
+(0, 5E-3)
+(80, 3.78)
.ENDS VCVS_LIMIT_2 



*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_4  VC+ VC- IOUT+ IOUT-
*              
.PARAM GAIN = 100U
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS VCCS_LIMIT_4 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_5  VC+ VC- IOUT+ IOUT-
*              
.PARAM GAIN = .15
.PARAM INEG = -5
.PARAM IPOS= 6.88
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS VCCS_LIMIT_5 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_1  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E6
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_1 


.END
