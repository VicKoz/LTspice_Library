* TLC271M OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.03 ON 06/01/90 AT 08:17
* REV (N/A)      SUPPLY VOLTAGE: +/-5V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT TLC271M  1 2 3 4 5
*
  C1   11 12 6.62E-12
  C2    6  7 20.00E-12
  CPSR 85 86 79.6E-9
  DCM+ 81 82 DX
  DCM- 83 81 DX
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  ECMR 84 99 (2,99)  1
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  EPSR 85 0 POLY(1) (3,4) -244.8E-6  24.48E-6
  ENSE 89 2 POLY(1) (88,0) 1.1E-3  1
  FB 7 99 POLY(6) VB VC VE VLP VLN VPSR 0 33.77E6 -90E6 90E6 90E6 -90E6 33.7E6
  GA    6  0 11 12 54.66E-6
  GCM 0  6 10 99 2.181E-9
  GPSR 85 86 (85,86) 100E-6
  GRD1 60 11 (60,11) 5.467E-5
  GRD2 60 12 (60,12) 5.467E-5
  HLIM 90  0 VLIM 1K
  HCMR 80 1 POLY(2) VCM+ VCM- 0 1E2 1E2
  IRP 3 4 131.8E-6
  ISS   3 10 DC 11.20E-6
  IIO 2 0 .1E-12
  I1 88 0 1E-21
  J1   11  89 10 JX
  J2   12  80 10 JX
  R2    6  9 100.0E3
  RCM 84 81 1K
  RN1 88 0 45E3
  RO1   8  5 75
  RO2   7 99 75
  RSS  10 99 17.86E6
  VAD  60 4 -.4
  VCM+ 82 99 3.65
  VCM- 83 99 -4.75
  VB    9  0 DC 0
  VC    3 53 DC 2
  VE   54  4 DC .7
  VLIM  7  8 DC 0
  VLP  91  0 DC 25
  VLN   0 92 DC 25
  VPSR 0 86 DC 0
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=350.0E-15 BETA=533.6E-6 VTO=-.033 KF=9.0E-17)
.ENDS