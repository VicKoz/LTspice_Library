* ADG633 ����������� ������� �� ������ ������� ADG659 � ADG1236
* �������� ���� ���� SPDT �� ������ ADG659.cir
* �������� ����������
* ���������� ������� ������� �� ������ ADG1236.cir
* �������� ����, ���������� ������ ������� 
* Developed by: ViKo 
* Revision History: 2017.01

****************
* Connections
*	1 = SA
*	2 = SB
*	3 = D
*	4 = VIN (Low On SA-D, High On SB-D)
*	5 = VDD
*	6 = GND
*	7 = VSS
*	8 = /EN (Low On)
****************
.SUBCKT ADG633  1 2 3 4 5 6 7 8
X1 1 3 4 5 6 7 8 LOWONSWITCH
X2 2 3 4 5 6 7 8 HIGHONSWITCH
RL1 5 6 5000MEG
RL2 7 6 5000MEG
CEN 8 6 2p
CIN 4 6 2p
DENA 8 5 DY
DENB 7 8 DY
DINA 4 5 DY
DINB 7 4 DY
CAB 1 2 0.15p

*MODELS USED
.MODEL DY D(IS=1E-14 N=0.04 RS=30)
.ENDS

****************
* Logic High On Switch
* Connections
*	101 = S
*	102 = D
*	103 = VIN
*	104 = VDD 
*	105 = GND
*	106 = VSS
*	107 = /EN
*****************
.SUBCKT HIGHONSWITCH  101 102 103 104 105 106 107
X1 103 104 105 108 BUFF
X2 108 109 104 106 105 VSENSE
X3 109 110 107 105 ENABLE
X4 110 105 111 ENABLEDELAY
X5 101 102 111 104 105 106 SWITCH

*MODELS USED
.ENDS

****************
* Logic Low On Switch
* Connections
*	101 = S
*	102 = D
*	103 = VIN
*	104 = VDD
*	105 = GND
*	106 = VSS
*	107 = /EN
****************
.SUBCKT LOWONSWITCH  101 102 103 104 105 106 107
X1 103 104 105 108 NOTGATE
X2 108 109 104 106 105 VSENSE
X3 109 110 107 105 ENABLE
X4 110 105 111 ENABLEDELAY
X5 101 102 111 104 105 106 SWITCH

*MODELS USED
.ENDS

****************
* Switch
* Connections
*	201 = S
*	202 = D
*	203 = VIN
*	204 = VDD 
*	205 = GND
*	206 = VSS
*****************
.SUBCKT SWITCH  201 202 203 204 205 206

*ANALOG SWITCH
EBuffer 214 205 202 205 1
S1 210 202 203 205 SMOD1
Vo2 214 219 0
EVDD 219 220 204 205 1
SN 210 209 205 220 SMOD7
Vo1 205 218 0
EVSS 217 218 206 205 1
SP 210 208 214 217 SMOD8 
Xn 215 209 214 205 204 206 VCRN
Xp 207 208 214 205 204 206 VCRP
RS1 201 207 1
RS2 201 215 1

DS1 201 204 DX 
DS2 206 201 DX
DD1 202 204 DX
DD2 206 202 DX

*ON OFF ISOLATION
CSD 201 202 0.201p
 
*BANDWIDTH 
CSB 201 206 2.1p
CDB 202 204 2.1p

*CHARGE INJECTION
CGS 201 203 0.167p
CGD 202 203 0.167p

*MODELS USED
.MODEL SMOD1 VSWITCH(RON=1 ROFF=7E11 VON=2.0 VOFF=0.8)
.MODEL SMOD7 VSWITCH(RON=1E-3 ROFF=1E11 VON=0.81 VOFF=0.79)
.MODEL SMOD8 VSWITCH(RON=1E-3 ROFF=1E11 VON=1.21 VOFF=1.19)
.MODEL DX D(IS=1E-12 N=0.04 RS=120)
.ENDS

*****************
* BUFF LOGIC
* Connections
*	201 = INPUT
*	202 = VDD
*	203 = GND
*	204 = OUTPUT
*****************
.SUBCKT BUFF 201 202 203 204
SBUFF 205 203 201 203 SMOD2
RBUFF 205 202 5G
EBUFFER 204 203 205 203 1

*MODELS USED
.MODEL SMOD2 VSWITCH(RON=1E-3 ROFF=1E11 VON=0.8 VOFF=2.0)
.ENDS

*****************
* NOT LOGIC
* Connections
*	201 = INPUT
*	202 = VDD
*	203 = GND
*	204 = OUTPUT
*****************
.SUBCKT NOTGATE 201 202 203 204
SNOT 205 203 201 203 SMOD2
RNOT 205 202 5G
EBUFFER 204 203 205 203 1

*MODELS USED
.MODEL SMOD2 VSWITCH(RON=1E-3 ROFF=1E11 VON=2.0 VOFF=0.8)
.ENDS

*****************
* ENABLE DELAY
* Connections
*	301 = INPUT
*	302 = COM
*	303 = OUTPUT
*****************
.SUBCKT ENABLEDELAY 301 302 303
EENBUFFER 304 302 301 302 1
RFEN 304 306 45k
CFEN 306 302 5p
DBREAKEN 306 305 DZ
RBEN 305 304 17k
EENBUFFEROUT 303 302 306 302 1 

*MODELS USED
.MODEL DZ D(IS=1E-14 N=0.04)
.ENDS

*****************
* Enable ON/OFF 
* Connections
*	501 = INPUT
*	502 = OUTPUT
*	503 = VIN
*	504 = GND
*****************
.SUBCKT ENABLE 501 502 503 504 
SENABLE 501 505 503 504 SMOD2
RD0 505 504 5G
EBUFFER 502 504 505 504 1

*MODELS USED
.MODEL SMOD2 VSWITCH(RON=1E-3 ROFF=1E11 VON=0.8 VOFF=2.0)
.ENDS

*****************
* OPERATING VOLTAGE 
* Connections
*	601 = INPUT
*	602 = OUTPUT
*	603 = VDD
*	604 = VSS
*	605 = GND
*****************
.SUBCKT VSENSE 601 602 603 604 605
SD1 601 606 603 605 SMOD3
SD2 606 607 603 605 SMOD4
SD3 607 608 605 604 SMOD5
SD4 608 609 605 604 SMOD6
SD5 609 602 603 604 SMOD7
RD0 602 605 5G

*MODELS USED
.MODEL SMOD3 VSWITCH(RON=1E-3 ROFF=1E11 VON=2 VOFF=1.9)
.MODEL SMOD4 VSWITCH(RON=1E-3 ROFF=1E11 VON=12 VOFF=12.1)
.MODEL SMOD5 VSWITCH(RON=1E-3 ROFF=1E11 VON=0 VOFF=-0.1)
.MODEL SMOD6 VSWITCH(RON=1E-3 ROFF=1E11 VON=6 VOFF=6.1)
.MODEL SMOD7 VSWITCH(RON=1E-3 ROFF=1E11 VON=12 VOFF=12.1)
.ENDS

*****************
* Voltage Controlled Resistance n-channel
* Connections
*	701 = R+
*	702 = R-
*	704 = V+
*	705 = V-
*	707 = VDD
*	711 = VSS
*****************
.SUBCKT VCRN 701 702 704 705 707 711
vtn 708 0 0.8
ERES 701 703 VALUE={285*V(706,0)*(1/(V(707,0)-V(704,705)-V(708,0)))}
VSENSE 703 702 0
FCOPY 0 706 VSENSE 1
RRES 706 0 1
.ENDS

*****************
* Voltage Controlled Resistance p-channel
* Connections
*	701 = R+
*	702 = R-
*	704 = V+
*	705 = V-
*	707 = VDD
*	711 = VSS
*****************
.SUBCKT VCRP 701 702 704 705 707 711
vtp 708 0 1.2
ERES 701 703 VALUE={246*V(706,0)*(1/(V(704,705)-V(711,0)-V(708,0)))}
VSENSE 703 702 0
FCOPY 0 706 VSENSE 1
RRES 706 0 1
.ENDS




